/*
 *  Control logic
 */
`default_nettype none
module control (ALU_Op, ALU_Src, instr);

    output wire ALU_Op, ALU_Src;

    input [15:0] instr;


    always @ (*) begin

    end


endmodule
`default_nettype wire
